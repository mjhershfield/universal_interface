module usb
    ();

endmodule
