module arbiter
    ();
    
endmodule
